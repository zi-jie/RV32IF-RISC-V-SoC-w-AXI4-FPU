`include "CPU_wrapper.sv"
`include "../src/AXI/AXI.sv"
`include "SRAM_wrapper.sv" // S1, S2
`include "ROM_wrapper.sv"  // S0
`include "DMA_wrapper.sv"  // S3
`include "WDT_wrapper.sv"  // S4
`include "DRAM_wrapper.sv" // S5

module top (
	input clk,
	input rst,
	input clk2,
	input rst2,
	// connect with ROM
	input [31:0] ROM_out,
	output logic ROM_read,
	output logic ROM_enable,
	output logic [11:0] ROM_address,
	// connect with DRAM
	input [31:0] DRAM_Q,
	input DRAM_valid,
	output logic DRAM_CSn,
	output logic [3:0] DRAM_WEn,
	output logic DRAM_RASn,
	output logic DRAM_CASn,
	output logic [10:0] DRAM_A,
	output logic [31:0] DRAM_D
);

logic DMA_interrupt;
logic WDT_interrupt;

/* Master */
// Master 1: AW
logic [`AXI_ID_BITS-1:0]    AWID_M1;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_M1;
logic [`AXI_LEN_BITS-1:0]   AWLEN_M1;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_M1;
logic [1:0]                 AWBURST_M1;
logic                       AWVALID_M1;
logic                       AWREADY_M1;
// Master 1: W
logic [`AXI_DATA_BITS-1:0]  WDATA_M1;
logic [`AXI_STRB_BITS-1:0]  WSTRB_M1;
logic                       WLAST_M1;
logic                       WVALID_M1;
logic                       WREADY_M1;
logic [`AXI_ID_BITS-1:0]    BID_M1;
logic [1:0]                 BRESP_M1;
logic                       BVALID_M1;
logic                       BREADY_M1;
// Master 0: AR
logic [`AXI_ID_BITS-1:0]    ARID_M0;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_M0;
logic [`AXI_LEN_BITS-1:0]   ARLEN_M0;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_M0;
logic [1:0]                 ARBURST_M0;
logic                       ARVALID_M0;
logic                       ARREADY_M0;
// Master 0: R
logic [`AXI_ID_BITS-1:0]    RID_M0;
logic [`AXI_DATA_BITS-1:0]  RDATA_M0;
logic [1:0]                 RRESP_M0;
logic                       RLAST_M0;
logic                       RVALID_M0;
logic                       RREADY_M0;
// Master 1: AR
logic [`AXI_ID_BITS-1:0]    ARID_M1;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_M1;
logic [`AXI_LEN_BITS-1:0]   ARLEN_M1;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_M1;
logic [1:0]                 ARBURST_M1;
logic                       ARVALID_M1;
logic                       ARREADY_M1;
// Master 1: R
logic [`AXI_ID_BITS-1:0]    RID_M1;
logic [`AXI_DATA_BITS-1:0]  RDATA_M1;
logic [1:0]                 RRESP_M1;
logic                       RLAST_M1;
logic                       RVALID_M1;
logic                       RREADY_M1;

/* Master 2 */
// Master 2 (DMA): AW
logic [`AXI_ID_BITS-1:0]    AWID_M2;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_M2;
logic [`AXI_LEN_BITS-1:0]   AWLEN_M2;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_M2;
logic [1:0]                 AWBURST_M2;
logic                       AWVALID_M2;
logic                       AWREADY_M2;
// Master 2 (DMA): W
logic [`AXI_DATA_BITS-1:0]  WDATA_M2;
logic [`AXI_STRB_BITS-1:0]  WSTRB_M2;
logic                       WLAST_M2;
logic                       WVALID_M2;
logic                       WREADY_M2;
logic [`AXI_ID_BITS-1:0]    BID_M2;
logic [1:0]                 BRESP_M2;
logic                       BVALID_M2;
logic                       BREADY_M2;
// Master 2 (DMA): AR
logic [`AXI_ID_BITS-1:0]    ARID_M2;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_M2;
logic [`AXI_LEN_BITS-1:0]   ARLEN_M2;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_M2;
logic [1:0]                 ARBURST_M2;
logic                       ARVALID_M2;
logic                       ARREADY_M2;
// Master 2 (DMA): R
logic [`AXI_ID_BITS-1:0]    RID_M2;
logic [`AXI_DATA_BITS-1:0]  RDATA_M2;
logic [1:0]                 RRESP_M2;
logic                       RLAST_M2;
logic                       RVALID_M2;
logic                       RREADY_M2;

/* Slave */
// Slave 1: AW
logic [`AXI_IDS_BITS-1:0]   AWID_S1;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_S1;
logic [`AXI_LEN_BITS-1:0]   AWLEN_S1;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_S1;
logic [1:0]                 AWBURST_S1;
logic                       AWVALID_S1;
logic                       AWREADY_S1;
// Slave 1: W
logic [`AXI_DATA_BITS-1:0]  WDATA_S1;
logic [`AXI_STRB_BITS-1:0]  WSTRB_S1;
logic                       WLAST_S1;
logic                       WVALID_S1;
logic                       WREADY_S1;
// Slave 1: B
logic [`AXI_IDS_BITS-1:0]   BID_S1;
logic [1:0]                 BRESP_S1;
logic                       BVALID_S1;
logic                       BREADY_S1;
// Slave 2: AW
logic [`AXI_IDS_BITS-1:0]   AWID_S2;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_S2;
logic [`AXI_LEN_BITS-1:0]   AWLEN_S2;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_S2;
logic [1:0]                 AWBURST_S2;
logic                       AWVALID_S2;
logic                       AWREADY_S2;
// Slave 2: W   
logic [`AXI_DATA_BITS-1:0]  WDATA_S2;
logic [`AXI_STRB_BITS-1:0]  WSTRB_S2;
logic                       WLAST_S2;
logic                       WVALID_S2;
logic                       WREADY_S2;
// Slave 2: B
logic [`AXI_IDS_BITS-1:0]   BID_S2;
logic [1:0]                 BRESP_S2;
logic                       BVALID_S2;
logic                       BREADY_S2;
// Slave 1: AR
logic [`AXI_IDS_BITS-1:0]   ARID_S1;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_S1;
logic [`AXI_LEN_BITS-1:0]   ARLEN_S1;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_S1;
logic [1:0]                 ARBURST_S1;
logic                       ARVALID_S1;
logic                       ARREADY_S1;
// Slave 1: R
logic [`AXI_IDS_BITS-1:0]   RID_S1;
logic [`AXI_DATA_BITS-1:0]  RDATA_S1;
logic [1:0]                 RRESP_S1;
logic                       RLAST_S1;
logic                       RVALID_S1;
logic                       RREADY_S1;
// Slave 2: AR
logic [`AXI_IDS_BITS-1:0]   ARID_S2;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_S2;
logic [`AXI_LEN_BITS-1:0]   ARLEN_S2;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_S2;
logic [1:0]                 ARBURST_S2;
logic                       ARVALID_S2;
logic                       ARREADY_S2;
// Slave 2: R
logic [`AXI_IDS_BITS-1:0]   RID_S2;
logic [`AXI_DATA_BITS-1:0]  RDATA_S2;
logic [1:0]                 RRESP_S2;
logic                       RLAST_S2;
logic                       RVALID_S2;
logic                       RREADY_S2;

/* Slave 0 */
// Slave 0 (ROM): AR
logic [`AXI_IDS_BITS-1:0]   ARID_S0;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_S0;
logic [`AXI_LEN_BITS-1:0]   ARLEN_S0;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_S0;
logic [1:0]                 ARBURST_S0;
logic                       ARVALID_S0;
logic                       ARREADY_S0;
// Slave 0 (ROM): R
logic [`AXI_IDS_BITS-1:0]   RID_S0;
logic [`AXI_DATA_BITS-1:0]  RDATA_S0;
logic [1:0]                 RRESP_S0;
logic                       RLAST_S0;
logic                       RVALID_S0;
logic                       RREADY_S0;

/* Slave 3 */
// Slave 3 (DMA): AW
logic [`AXI_IDS_BITS-1:0]   AWID_S3;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_S3;
logic [`AXI_LEN_BITS-1:0]   AWLEN_S3;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_S3;
logic [1:0]                 AWBURST_S3;
logic                       AWVALID_S3;
logic                       AWREADY_S3;
// Slave 3 (DMA): W   
logic [`AXI_DATA_BITS-1:0]  WDATA_S3;
logic [`AXI_STRB_BITS-1:0]  WSTRB_S3;
logic                       WLAST_S3;
logic                       WVALID_S3;
logic                       WREADY_S3;
// Slave 3 (DMA): B
logic [`AXI_IDS_BITS-1:0]   BID_S3;
logic [1:0]                 BRESP_S3;
logic                       BVALID_S3;
logic                       BREADY_S3;

/* Slave 4: WDT */ 
// AW
logic [`AXI_IDS_BITS-1:0]   AWID_S4;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_S4;
logic [`AXI_LEN_BITS-1:0]   AWLEN_S4;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_S4;
logic [1:0]                 AWBURST_S4;
logic                       AWVALID_S4;
logic                       AWREADY_S4;
// W
logic [`AXI_DATA_BITS-1:0]  WDATA_S4;
logic [`AXI_STRB_BITS-1:0]  WSTRB_S4;
logic                       WLAST_S4;
logic                       WVALID_S4;
logic                       WREADY_S4;
// B
logic [`AXI_IDS_BITS-1:0]   BID_S4;
logic [1:0]                 BRESP_S4;
logic                       BVALID_S4;
logic                       BREADY_S4;
// AR
logic [`AXI_IDS_BITS-1:0]   ARID_S4;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_S4;
logic [`AXI_LEN_BITS-1:0]   ARLEN_S4;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_S4;
logic [1:0]                 ARBURST_S4;
logic                       ARVALID_S4;
logic                       ARREADY_S4;
// R
logic [`AXI_IDS_BITS-1:0]   RID_S4;
logic [`AXI_DATA_BITS-1:0]  RDATA_S4;
logic [1:0]                 RRESP_S4;
logic                       RLAST_S4;
logic                       RVALID_S4;
logic                       RREADY_S4;

/* Slave 5: DRAM */
// Slave 5 (DRAM): AW
logic [`AXI_IDS_BITS-1:0]   AWID_S5;
logic [`AXI_ADDR_BITS-1:0]  AWADDR_S5;
logic [`AXI_LEN_BITS-1:0]   AWLEN_S5;
logic [`AXI_SIZE_BITS-1:0]  AWSIZE_S5;
logic [1:0]                 AWBURST_S5;
logic                       AWVALID_S5;
logic                       AWREADY_S5;
// Slave 5 (DRAM): W   
logic [`AXI_DATA_BITS-1:0]  WDATA_S5;
logic [`AXI_STRB_BITS-1:0]  WSTRB_S5;
logic                       WLAST_S5;
logic                       WVALID_S5;
logic                       WREADY_S5;
// Slave 5 (DRAM): B
logic [`AXI_IDS_BITS-1:0]   BID_S5;
logic [1:0]                 BRESP_S5;
logic                       BVALID_S5;
logic                       BREADY_S5;
// Slave 5 (DRAM): AR
logic [`AXI_IDS_BITS-1:0]   ARID_S5;
logic [`AXI_ADDR_BITS-1:0]  ARADDR_S5;
logic [`AXI_LEN_BITS-1:0]   ARLEN_S5;
logic [`AXI_SIZE_BITS-1:0]  ARSIZE_S5;
logic [1:0]                 ARBURST_S5;
logic                       ARVALID_S5;
logic                       ARREADY_S5;
// Slave 5 (DRAM): R
logic [`AXI_IDS_BITS-1:0]   RID_S5;
logic [`AXI_DATA_BITS-1:0]  RDATA_S5;
logic [1:0]                 RRESP_S5;
logic                       RLAST_S5;
logic                       RVALID_S5;
logic                       RREADY_S5;

CPU_wrapper CPU_wrapper1(
	.ACLK(clk),
	.ARESETn(~rst),
	.DMA_interrupt(DMA_interrupt),
	// .WDT_interrupt(1'b0), //FIXME: 0 -> WDT_interrupt
	.WDT_interrupt(WDT_interrupt), 
	.AWID_M1(AWID_M1),
	.AWADDR_M1(AWADDR_M1),
	.AWLEN_M1(AWLEN_M1),
	.AWSIZE_M1(AWSIZE_M1),
	.AWBURST_M1(AWBURST_M1),
	.AWVALID_M1(AWVALID_M1),
	.AWREADY_M1(AWREADY_M1),		
	.WDATA_M1(WDATA_M1),     
	.WSTRB_M1(WSTRB_M1), 
	.WLAST_M1(WLAST_M1),
	.WVALID_M1(WVALID_M1),
	.WREADY_M1(WREADY_M1),
	.BID_M1(BID_M1),
	.BRESP_M1(BRESP_M1),
	.BVALID_M1(BVALID_M1),
	.BREADY_M1(BREADY_M1), 
	.ARID_M0(ARID_M0),
	.ARADDR_M0(ARADDR_M0),
	.ARLEN_M0(ARLEN_M0),
	.ARSIZE_M0(ARSIZE_M0),
	.ARBURST_M0(ARBURST_M0),
	.ARVALID_M0(ARVALID_M0),
	.ARREADY_M0(ARREADY_M0),
	.RID_M0(RID_M0),		
	.RDATA_M0(RDATA_M0),
	.RRESP_M0(RRESP_M0),
	.RLAST_M0(RLAST_M0),
	.RVALID_M0(RVALID_M0),
	.RREADY_M0(RREADY_M0),
	.ARID_M1(ARID_M1),
	.ARADDR_M1(ARADDR_M1),
	.ARLEN_M1(ARLEN_M1),
	.ARSIZE_M1(ARSIZE_M1),
	.ARBURST_M1(ARBURST_M1),
	.ARVALID_M1(ARVALID_M1),
	.ARREADY_M1(ARREADY_M1),
	.RID_M1(RID_M1),
	.RDATA_M1(RDATA_M1),
	.RRESP_M1(RRESP_M1),
	.RLAST_M1(RLAST_M1),
	.RVALID_M1(RVALID_M1),
	.RREADY_M1(RREADY_M1)    
);

//TODO: connect AXI
AXI AXI1(
	.ACLK(clk),
	.ARESETn(~rst),
	.AWID_M1(AWID_M1),
	.AWADDR_M1(AWADDR_M1),
	.AWLEN_M1(AWLEN_M1),
	.AWSIZE_M1(AWSIZE_M1),
	.AWBURST_M1(AWBURST_M1),
	.AWVALID_M1(AWVALID_M1),
	.AWREADY_M1(AWREADY_M1),
	.WDATA_M1(WDATA_M1),
	.WSTRB_M1(WSTRB_M1),
	.WLAST_M1(WLAST_M1),
	.WVALID_M1(WVALID_M1),
	.WREADY_M1(WREADY_M1),
	.BID_M1(BID_M1),
	.BRESP_M1(BRESP_M1),
	.BVALID_M1(BVALID_M1),
	.BREADY_M1(BREADY_M1),
	.AWID_M2(AWID_M2),
	.AWADDR_M2(AWADDR_M2),
	.AWLEN_M2(AWLEN_M2),
	.AWSIZE_M2(AWSIZE_M2),
	.AWBURST_M2(AWBURST_M2),
	.AWVALID_M2(AWVALID_M2),
	.AWREADY_M2(AWREADY_M2),
	.WDATA_M2(WDATA_M2),
	.WSTRB_M2(WSTRB_M2),
	.WLAST_M2(WLAST_M2),
	.WVALID_M2(WVALID_M2),
	.WREADY_M2(WREADY_M2),
	.BID_M2(BID_M2),
	.BRESP_M2(BRESP_M2),
	.BVALID_M2(BVALID_M2),
	.BREADY_M2(BREADY_M2),
	.ARID_M0(ARID_M0),
	.ARADDR_M0(ARADDR_M0),
	.ARLEN_M0(ARLEN_M0),
	.ARSIZE_M0(ARSIZE_M0),
	.ARBURST_M0(ARBURST_M0),
	.ARVALID_M0(ARVALID_M0),
	.ARREADY_M0(ARREADY_M0),
	.RID_M0(RID_M0),
	.RDATA_M0(RDATA_M0),
	.RRESP_M0(RRESP_M0),
	.RLAST_M0(RLAST_M0),
	.RVALID_M0(RVALID_M0),
	.RREADY_M0(RREADY_M0),
	.ARID_M1(ARID_M1),
	.ARADDR_M1(ARADDR_M1),
	.ARLEN_M1(ARLEN_M1),
	.ARSIZE_M1(ARSIZE_M1),
	.ARBURST_M1(ARBURST_M1),
	.ARVALID_M1(ARVALID_M1),
	.ARREADY_M1(ARREADY_M1),
	.RID_M1(RID_M1),
	.RDATA_M1(RDATA_M1),
	.RRESP_M1(RRESP_M1),
	.RLAST_M1(RLAST_M1),
	.RVALID_M1(RVALID_M1),
	.RREADY_M1(RREADY_M1),
	.ARID_M2(ARID_M2),
	.ARADDR_M2(ARADDR_M2),
	.ARLEN_M2(ARLEN_M2),
	.ARSIZE_M2(ARSIZE_M2),
	.ARBURST_M2(ARBURST_M2),
	.ARVALID_M2(ARVALID_M2),
	.ARREADY_M2(ARREADY_M2),
	.RID_M2(RID_M2),
	.RDATA_M2(RDATA_M2),
	.RRESP_M2(RRESP_M2),
	.RLAST_M2(RLAST_M2),
	.RVALID_M2(RVALID_M2),
	.RREADY_M2(RREADY_M2),
	.AWID_S1(AWID_S1),
	.AWADDR_S1(AWADDR_S1),
	.AWLEN_S1(AWLEN_S1),
	.AWSIZE_S1(AWSIZE_S1),
	.AWBURST_S1(AWBURST_S1),
	.AWVALID_S1(AWVALID_S1),
	.AWREADY_S1(AWREADY_S1),
	.WDATA_S1(WDATA_S1),
	.WSTRB_S1(WSTRB_S1),
	.WLAST_S1(WLAST_S1),
	.WVALID_S1(WVALID_S1),
	.WREADY_S1(WREADY_S1),
	.BID_S1(BID_S1),
	.BRESP_S1(BRESP_S1),
	.BVALID_S1(BVALID_S1),
	.BREADY_S1(BREADY_S1),
	.AWID_S2(AWID_S2),
	.AWADDR_S2(AWADDR_S2),
	.AWLEN_S2(AWLEN_S2),
	.AWSIZE_S2(AWSIZE_S2),
	.AWBURST_S2(AWBURST_S2),
	.AWVALID_S2(AWVALID_S2),
	.AWREADY_S2(AWREADY_S2),
	.WDATA_S2(WDATA_S2),
	.WSTRB_S2(WSTRB_S2),
	.WLAST_S2(WLAST_S2),
	.WVALID_S2(WVALID_S2),
	.WREADY_S2(WREADY_S2),
	.BID_S2(BID_S2),
	.BRESP_S2(BRESP_S2),
	.BVALID_S2(BVALID_S2),
	.BREADY_S2(BREADY_S2),
	.AWID_S3(AWID_S3),
	.AWADDR_S3(AWADDR_S3),
	.AWLEN_S3(AWLEN_S3),
	.AWSIZE_S3(AWSIZE_S3),
	.AWBURST_S3(AWBURST_S3),
	.AWVALID_S3(AWVALID_S3),
	.AWREADY_S3(AWREADY_S3),
	.WDATA_S3(WDATA_S3),
	.WSTRB_S3(WSTRB_S3),
	.WLAST_S3(WLAST_S3),
	.WVALID_S3(WVALID_S3),
	.WREADY_S3(WREADY_S3),
	.BID_S3(BID_S3),
	.BRESP_S3(BRESP_S3),
	.BVALID_S3(BVALID_S3),
	.BREADY_S3(BREADY_S3),
	.AWID_S4(AWID_S4),
	.AWADDR_S4(AWADDR_S4),
	.AWLEN_S4(AWLEN_S4),
	.AWSIZE_S4(AWSIZE_S4),
	.AWBURST_S4(AWBURST_S4),
	.AWVALID_S4(AWVALID_S4),
	.AWREADY_S4(AWREADY_S4),
	.WDATA_S4(WDATA_S4),
	.WSTRB_S4(WSTRB_S4),
	.WLAST_S4(WLAST_S4),
	.WVALID_S4(WVALID_S4),
	.WREADY_S4(WREADY_S4),
	.BID_S4(BID_S4),
	.BRESP_S4(BRESP_S4),
	.BVALID_S4(BVALID_S4),
	.BREADY_S4(BREADY_S4),
	.AWID_S5(AWID_S5),
	.AWADDR_S5(AWADDR_S5),
	.AWLEN_S5(AWLEN_S5),
	.AWSIZE_S5(AWSIZE_S5),
	.AWBURST_S5(AWBURST_S5),
	.AWVALID_S5(AWVALID_S5),
	.AWREADY_S5(AWREADY_S5),
	.WDATA_S5(WDATA_S5),
	.WSTRB_S5(WSTRB_S5),
	.WLAST_S5(WLAST_S5),
	.WVALID_S5(WVALID_S5),
	.WREADY_S5(WREADY_S5),
	.BID_S5(BID_S5),
	.BRESP_S5(BRESP_S5),
	.BVALID_S5(BVALID_S5),
	.BREADY_S5(BREADY_S5),
	.ARID_S0(ARID_S0),
	.ARADDR_S0(ARADDR_S0),
	.ARLEN_S0(ARLEN_S0),
	.ARSIZE_S0(ARSIZE_S0),
	.ARBURST_S0(ARBURST_S0),
	.ARVALID_S0(ARVALID_S0),
	.ARREADY_S0(ARREADY_S0),
	.RID_S0(RID_S0),
	.RDATA_S0(RDATA_S0),
	.RRESP_S0(RRESP_S0),
	.RLAST_S0(RLAST_S0),
	.RVALID_S0(RVALID_S0),
	.RREADY_S0(RREADY_S0),
	.ARID_S1(ARID_S1),
	.ARADDR_S1(ARADDR_S1),
	.ARLEN_S1(ARLEN_S1),
	.ARSIZE_S1(ARSIZE_S1),
	.ARBURST_S1(ARBURST_S1),
	.ARVALID_S1(ARVALID_S1),
	.ARREADY_S1(ARREADY_S1),
	.RID_S1(RID_S1),
	.RDATA_S1(RDATA_S1),
	.RRESP_S1(RRESP_S1),
	.RLAST_S1(RLAST_S1),
	.RVALID_S1(RVALID_S1),
	.RREADY_S1(RREADY_S1),
	.ARID_S2(ARID_S2),
	.ARADDR_S2(ARADDR_S2),
	.ARLEN_S2(ARLEN_S2),
	.ARSIZE_S2(ARSIZE_S2),
	.ARBURST_S2(ARBURST_S2),
	.ARVALID_S2(ARVALID_S2),
	.ARREADY_S2(ARREADY_S2),
	.RID_S2(RID_S2),
	.RDATA_S2(RDATA_S2),
	.RRESP_S2(RRESP_S2),
	.RLAST_S2(RLAST_S2),
	.RVALID_S2(RVALID_S2),
	.RREADY_S2(RREADY_S2),
	.ARID_S4(ARID_S4),
	.ARADDR_S4(ARADDR_S4),
	.ARLEN_S4(ARLEN_S4),
	.ARSIZE_S4(ARSIZE_S4),
	.ARBURST_S4(ARBURST_S4),
	.ARVALID_S4(ARVALID_S4),
	.ARREADY_S4(ARREADY_S4),
	.RID_S4(RID_S4),
	.RDATA_S4(RDATA_S4),
	.RRESP_S4(RRESP_S4),
	.RLAST_S4(RLAST_S4),
	.RVALID_S4(RVALID_S4),
	.RREADY_S4(RREADY_S4),
	.ARID_S5(ARID_S5),
	.ARADDR_S5(ARADDR_S5),
	.ARLEN_S5(ARLEN_S5),
	.ARSIZE_S5(ARSIZE_S5),
	.ARBURST_S5(ARBURST_S5),
	.ARVALID_S5(ARVALID_S5),
	.ARREADY_S5(ARREADY_S5),
	.RID_S5(RID_S5),
	.RDATA_S5(RDATA_S5),
	.RRESP_S5(RRESP_S5),
	.RLAST_S5(RLAST_S5),
	.RVALID_S5(RVALID_S5),
	.RREADY_S5(RREADY_S5)
);

// Slave 0: ROM (only read)
ROM_wrapper ROM1(
    .ACLK(clk),
    .ARESETn(~rst),
    .ARID_S0(ARID_S0),     
    .ARADDR_S0(ARADDR_S0),       
    .ARLEN_S0(ARLEN_S0),       
    .ARSIZE_S0(ARSIZE_S0),       
    .ARBURST_S0(ARBURST_S0),      
    .ARVALID_S0(ARVALID_S0),      
    .ARREADY_S0(ARREADY_S0),      
    .RID_S0(RID_S0),
    .RDATA_S0(RDATA_S0),       
    .RRESP_S0(RRESP_S0),       
    .RLAST_S0(RLAST_S0),       
    .RVALID_S0(RVALID_S0),       
    .RREADY_S0(RREADY_S0),
    .ROM_out(ROM_out),
    .ROM_read(ROM_read),
    .ROM_enable(ROM_enable),
    .ROM_address(ROM_address)
);

// Slave 1
SRAM_wrapper IM1(
	.ACLK(clk),
	.ARESETn(~rst),
	.AWID_S(AWID_S1),
	.AWADDR_S(AWADDR_S1),    
	.AWLEN_S(AWLEN_S1),       
	.AWSIZE_S(AWSIZE_S1),       
	.AWBURST_S(AWBURST_S1),    
	.AWVALID_S(AWVALID_S1),
	.AWREADY_S(AWREADY_S1),    
	.WDATA_S(WDATA_S1),
	.WSTRB_S(WSTRB_S1),       
	.WLAST_S(WLAST_S1),       
	.WVALID_S(WVALID_S1),      
	.WREADY_S(WREADY_S1),      
	.BID_S(BID_S1),
	.BRESP_S(BRESP_S1),       
	.BVALID_S(BVALID_S1),       
	.BREADY_S(BREADY_S1),       
	.ARID_S(ARID_S1),     
	.ARADDR_S(ARADDR_S1),       
	.ARLEN_S(ARLEN_S1),       
	.ARSIZE_S(ARSIZE_S1),       
	.ARBURST_S(ARBURST_S1),      
	.ARVALID_S(ARVALID_S1),      
	.ARREADY_S(ARREADY_S1),      
	.RID_S(RID_S1),
	.RDATA_S(RDATA_S1),       
	.RRESP_S(RRESP_S1),       
	.RLAST_S(RLAST_S1),       
	.RVALID_S(RVALID_S1),       
	.RREADY_S(RREADY_S1)     
);

// Slave 2
SRAM_wrapper DM1(
	.ACLK(clk),
	.ARESETn(~rst),
	.AWID_S(AWID_S2),
	.AWADDR_S(AWADDR_S2),    
	.AWLEN_S(AWLEN_S2),       
	.AWSIZE_S(AWSIZE_S2),       
	.AWBURST_S(AWBURST_S2),    
	.AWVALID_S(AWVALID_S2),
	.AWREADY_S(AWREADY_S2),    
	.WDATA_S(WDATA_S2),
	.WSTRB_S(WSTRB_S2),       
	.WLAST_S(WLAST_S2),       
	.WVALID_S(WVALID_S2),      
	.WREADY_S(WREADY_S2),      
	.BID_S(BID_S2),
	.BRESP_S(BRESP_S2),       
	.BVALID_S(BVALID_S2),       
	.BREADY_S(BREADY_S2),       
	.ARID_S(ARID_S2),     
	.ARADDR_S(ARADDR_S2),       
	.ARLEN_S(ARLEN_S2),       
	.ARSIZE_S(ARSIZE_S2),       
	.ARBURST_S(ARBURST_S2),      
	.ARVALID_S(ARVALID_S2),      
	.ARREADY_S(ARREADY_S2),      
	.RID_S(RID_S2),
	.RDATA_S(RDATA_S2),       
	.RRESP_S(RRESP_S2),       
	.RLAST_S(RLAST_S2),       
	.RVALID_S(RVALID_S2),       
	.RREADY_S(RREADY_S2)   
);

// Slave 3: DMA (only write); Master 2
DMA_wrapper DMA1(
    .ACLK(clk),
    .ARESETn(~rst),
    .AWID_S3(AWID_S3), // Slave 3: only write channel
    .AWADDR_S3(AWADDR_S3),    
    .AWLEN_S3(AWLEN_S3),       
    .AWSIZE_S3(AWSIZE_S3),       
    .AWBURST_S3(AWBURST_S3),    
    .AWVALID_S3(AWVALID_S3),
    .AWREADY_S3(AWREADY_S3),    
    .WDATA_S3(WDATA_S3),
    .WSTRB_S3(WSTRB_S3),       
    .WLAST_S3(WLAST_S3),       
    .WVALID_S3(WVALID_S3),      
    .WREADY_S3(WREADY_S3),      
    .BID_S3(BID_S3),
    .BRESP_S3(BRESP_S3),       
    .BVALID_S3(BVALID_S3),       
    .BREADY_S3(BREADY_S3),
    .AWID_M2(AWID_M2),
    .AWADDR_M2(AWADDR_M2),
    .AWLEN_M2(AWLEN_M2),
    .AWSIZE_M2(AWSIZE_M2),
    .AWBURST_M2(AWBURST_M2),
    .AWVALID_M2(AWVALID_M2),
    .AWREADY_M2(AWREADY_M2),		
    .WDATA_M2(WDATA_M2),     
    .WSTRB_M2(WSTRB_M2), 
    .WLAST_M2(WLAST_M2),
    .WVALID_M2(WVALID_M2),
    .WREADY_M2(WREADY_M2),
    .BID_M2(BID_M2),
    .BRESP_M2(BRESP_M2),
    .BVALID_M2(BVALID_M2),
    .BREADY_M2(BREADY_M2), 
    .ARID_M2(ARID_M2),
    .ARADDR_M2(ARADDR_M2),
    .ARLEN_M2(ARLEN_M2),
    .ARSIZE_M2(ARSIZE_M2),
    .ARBURST_M2(ARBURST_M2),
    .ARVALID_M2(ARVALID_M2),
    .ARREADY_M2(ARREADY_M2),
    .RID_M2(RID_M2),		
    .RDATA_M2(RDATA_M2),
    .RRESP_M2(RRESP_M2),
    .RLAST_M2(RLAST_M2),
    .RVALID_M2(RVALID_M2),
    .RREADY_M2(RREADY_M2),
    .DMA_interrupt(DMA_interrupt) //TODO: connect with CPU
);

// Slave 4: WDT
WDT_wrapper WDT_wrapper1(
	.ACLK(clk),
	.ARESETn(~rst),
	.AWID_S(AWID_S4),
	.AWADDR_S(AWADDR_S4),    
	.AWLEN_S(AWLEN_S4),       
	.AWSIZE_S(AWSIZE_S4),       
	.AWBURST_S(AWBURST_S4),    
	.AWVALID_S(AWVALID_S4),
	.AWREADY_S(AWREADY_S4),    
	.WDATA_S(WDATA_S4),
	.WSTRB_S(WSTRB_S4),       
	.WLAST_S(WLAST_S4),       
	.WVALID_S(WVALID_S4),      
	.WREADY_S(WREADY_S4),      
	.BID_S(BID_S4),
	.BRESP_S(BRESP_S4),       
	.BVALID_S(BVALID_S4),       
	.BREADY_S(BREADY_S4),       
	.ARID_S(ARID_S4),     
	.ARADDR_S(ARADDR_S4),       
	.ARLEN_S(ARLEN_S4),       
	.ARSIZE_S(ARSIZE_S4),       
	.ARBURST_S(ARBURST_S4),      
	.ARVALID_S(ARVALID_S4),      
	.ARREADY_S(ARREADY_S4),      
	.RID_S(RID_S4),
	.RDATA_S(RDATA_S4),       
	.RRESP_S(RRESP_S4),       
	.RLAST_S(RLAST_S4),       
	.RVALID_S(RVALID_S4),       
	.RREADY_S(RREADY_S4),
	.clk2(clk2),
	.rst2(rst2),
	.WDT_interrupt(WDT_interrupt) //TODO: connect with CPU FIXME    
);

// Slave 5: DRAM
DRAM_wrapper DRAM1(
    .ACLK(clk),
    .ARESETn(~rst),
    .AWID_S5(AWID_S5),
    .AWADDR_S5(AWADDR_S5),    
    .AWLEN_S5(AWLEN_S5),       
    .AWSIZE_S5(AWSIZE_S5),       
    .AWBURST_S5(AWBURST_S5),    
    .AWVALID_S5(AWVALID_S5),
    .AWREADY_S5(AWREADY_S5),    
    .WDATA_S5(WDATA_S5),
    .WSTRB_S5(WSTRB_S5),       
    .WLAST_S5(WLAST_S5),       
    .WVALID_S5(WVALID_S5),      
    .WREADY_S5(WREADY_S5),      
    .BID_S5(BID_S5),
    .BRESP_S5(BRESP_S5),       
    .BVALID_S5(BVALID_S5),       
    .BREADY_S5(BREADY_S5),
    .ARID_S5(ARID_S5),     
    .ARADDR_S5(ARADDR_S5),       
    .ARLEN_S5(ARLEN_S5),       
    .ARSIZE_S5(ARSIZE_S5),       
    .ARBURST_S5(ARBURST_S5),      
    .ARVALID_S5(ARVALID_S5),      
    .ARREADY_S5(ARREADY_S5),      
    .RID_S5(RID_S5),
    .RDATA_S5(RDATA_S5),       
    .RRESP_S5(RRESP_S5),       
    .RLAST_S5(RLAST_S5),       
    .RVALID_S5(RVALID_S5),       
    .RREADY_S5(RREADY_S5),
    .DRAM_Q(DRAM_Q),
    .DRAM_valid(DRAM_valid),
    .DRAM_CSn(DRAM_CSn),
    .DRAM_WEn(DRAM_WEn),
    .DRAM_RASn(DRAM_RASn),
    .DRAM_CASn(DRAM_CASn),
    .DRAM_A(DRAM_A),
    .DRAM_D(DRAM_D)
);

endmodule