`define BANDWIDTH 32
`define MAC_NUM 9
`define PE_NUM 4
`define BYTE 8
`define HWORD 16
`define WORD 32
//mem config
`define IFM_MEM_SIZE 64
`define IFM_SIZE_BITS 6
`define WEIGHT_SIZE 3
`define OUT_BUF_SIZE 64
`define OUT_BUF_BITS 6
`define PE_BUF_SIZE 64 //PE_buffer 32*3 (*32)
